/***
 *                .-'''-.                              
 *               '   _    \                            
 *             /   /` '.   \    .        .--.          
 *            .   |     \  '  .'|        |__|          
 *    .-,.--. |   '      |  '<  |        .--.     .|   
 *    |  .-. |\    \     / /  | |        |  |   .' |_  
 *    | |  | | `.   ` ..' /   | | .'''-. |  | .'     | 
 *    | |  | |    '-...-'`    | |/.'''. \|  |'--.  .-' 
 *    | |  '-                 |  /    | ||  |   |  |   
 *    | |                     | |     | ||__|   |  |   
 *    | |                     | |     | |       |  '.' 
 *    |_|                     | '.    | '.      |   /  
 *                            '---'   '---'     `'-'   
 *
 *
 *	design: 	floating point (IEEE 754) multiplier without clk or reset, works with limited inputs
 *	date:		12.02.2018
 *	version:	1.0
 *
 */

// http://www.rfwireless-world.com/Tutorials/floating-point-tutorial.html
// http://www.ecs.umass.edu/ece/koren/arith/simulator/FPMul/
// http://weitz.de/ieee/

 module fpm #(parameter size = 32 )
 	(input logic [size-1 : 0] a, [size-1 : 0] b,
 	output logic [size-1 : 0] m
 	);

11001100110011001100110
11001100110011001100110

endmodule