// FPU